// Code for wire and logic 


module wire_logic;

wire a;
logic b;
reg c;

assign c=1;

assign a=1;
assign a=0;

initial
begin
	b=0;
end	

initial
begin
	b=1;
end
endmodule
