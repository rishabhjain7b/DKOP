// Code for understanding Interfaces with HA

interface ha_if;