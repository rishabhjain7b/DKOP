// Code interfacing 