// Code for testing type casting, size casting and  sign casting

module testcasting;