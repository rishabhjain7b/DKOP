// Code for testing ref keyword