// Code for assign in always

module test3;

reg a;

initial
begin
	assign a=1'b1;
	$display(a);
end
endmodule


