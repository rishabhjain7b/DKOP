// testbench of fork join

module fork_join_tb;
